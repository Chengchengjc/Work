`timescale 1ns/1ns
module Shifter( dataA, dataB, Signal, dataOut ) ;
input [31:0] dataA ;
input [31:0] dataB ;
input [5:0] Signal ;
output [31:0] dataOut ;

wire padding;
wire [31:0] temp, temp2, temp3, temp4, temp5 ;

assign padding = 1'b0;
parameter SRL = 6'b000010 ;

MUX2_1 m1 (.out(temp[0]), .in0(dataA[0]), .in1(dataA[1]), .sel(dataB[0])) ;
MUX2_1 m2 (.out(temp[1]), .in0(dataA[1]), .in1(dataA[2]), .sel(dataB[0])) ;
MUX2_1 m3 (.out(temp[2]), .in0(dataA[2]), .in1(dataA[3]), .sel(dataB[0])) ;
MUX2_1 m4 (.out(temp[3]), .in0(dataA[3]), .in1(dataA[4]), .sel(dataB[0])) ;
MUX2_1 m5 (.out(temp[4]), .in0(dataA[4]), .in1(dataA[5]), .sel(dataB[0])) ;
MUX2_1 m6 (.out(temp[5]), .in0(dataA[5]), .in1(dataA[6]), .sel(dataB[0])) ;
MUX2_1 m7 (.out(temp[6]), .in0(dataA[6]), .in1(dataA[7]), .sel(dataB[0])) ;
MUX2_1 m8 (.out(temp[7]), .in0(dataA[7]), .in1(dataA[8]), .sel(dataB[0])) ;
MUX2_1 m9 (.out(temp[8]), .in0(dataA[8]), .in1(dataA[9]), .sel(dataB[0])) ;
MUX2_1 m10 (.out(temp[9]), .in0(dataA[9]), .in1(dataA[10]), .sel(dataB[0])) ;
MUX2_1 m11 (.out(temp[10]), .in0(dataA[10]), .in1(dataA[11]), .sel(dataB[0])) ;
MUX2_1 m12 (.out(temp[11]), .in0(dataA[11]), .in1(dataA[12]), .sel(dataB[0])) ;
MUX2_1 m13 (.out(temp[12]), .in0(dataA[12]), .in1(dataA[13]), .sel(dataB[0])) ;
MUX2_1 m14 (.out(temp[13]), .in0(dataA[13]), .in1(dataA[14]), .sel(dataB[0])) ;
MUX2_1 m15 (.out(temp[14]), .in0(dataA[14]), .in1(dataA[15]), .sel(dataB[0])) ;
MUX2_1 m16 (.out(temp[15]), .in0(dataA[15]), .in1(dataA[16]), .sel(dataB[0])) ;
MUX2_1 m17 (.out(temp[16]), .in0(dataA[16]), .in1(dataA[17]), .sel(dataB[0])) ;
MUX2_1 m18 (.out(temp[17]), .in0(dataA[17]), .in1(dataA[18]), .sel(dataB[0])) ;
MUX2_1 m19 (.out(temp[18]), .in0(dataA[18]), .in1(dataA[19]), .sel(dataB[0])) ;
MUX2_1 m20 (.out(temp[19]), .in0(dataA[19]), .in1(dataA[20]), .sel(dataB[0])) ;
MUX2_1 m21 (.out(temp[20]), .in0(dataA[20]), .in1(dataA[21]), .sel(dataB[0])) ;
MUX2_1 m22 (.out(temp[21]), .in0(dataA[21]), .in1(dataA[22]), .sel(dataB[0])) ;
MUX2_1 m23 (.out(temp[22]), .in0(dataA[22]), .in1(dataA[23]), .sel(dataB[0])) ;
MUX2_1 m24 (.out(temp[23]), .in0(dataA[23]), .in1(dataA[24]), .sel(dataB[0])) ;
MUX2_1 m25 (.out(temp[24]), .in0(dataA[24]), .in1(dataA[25]), .sel(dataB[0])) ;
MUX2_1 m26 (.out(temp[25]), .in0(dataA[25]), .in1(dataA[26]), .sel(dataB[0])) ;
MUX2_1 m27 (.out(temp[26]), .in0(dataA[26]), .in1(dataA[27]), .sel(dataB[0])) ;
MUX2_1 m28 (.out(temp[27]), .in0(dataA[27]), .in1(dataA[28]), .sel(dataB[0])) ;
MUX2_1 m29 (.out(temp[28]), .in0(dataA[28]), .in1(dataA[29]), .sel(dataB[0])) ;
MUX2_1 m30 (.out(temp[29]), .in0(dataA[29]), .in1(dataA[30]), .sel(dataB[0])) ;
MUX2_1 m31 (.out(temp[30]), .in0(dataA[30]), .in1(dataA[31]), .sel(dataB[0])) ;
MUX2_1 m32 (.out(temp[31]), .in0(dataA[31]), .in1(padding), .sel(dataB[0])) ;

MUX2_1 m2_1 (.out(temp2[0]), .in0(temp[0]), .in1(temp[2]), .sel(dataB[1])) ;
MUX2_1 m2_2 (.out(temp2[1]), .in0(temp[1]), .in1(temp[3]), .sel(dataB[1])) ;
MUX2_1 m2_3 (.out(temp2[2]), .in0(temp[2]), .in1(temp[4]), .sel(dataB[1])) ;
MUX2_1 m2_4 (.out(temp2[3]), .in0(temp[3]), .in1(temp[5]), .sel(dataB[1])) ;
MUX2_1 m2_5 (.out(temp2[4]), .in0(temp[4]), .in1(temp[6]), .sel(dataB[1])) ;
MUX2_1 m2_6 (.out(temp2[5]), .in0(temp[5]), .in1(temp[7]), .sel(dataB[1])) ;
MUX2_1 m2_7 (.out(temp2[6]), .in0(temp[6]), .in1(temp[8]), .sel(dataB[1])) ;
MUX2_1 m2_8 (.out(temp2[7]), .in0(temp[7]), .in1(temp[9]), .sel(dataB[1])) ;
MUX2_1 m2_9 (.out(temp2[8]), .in0(temp[8]), .in1(temp[10]), .sel(dataB[1])) ;
MUX2_1 m2_10 (.out(temp2[9]), .in0(temp[9]), .in1(temp[11]), .sel(dataB[1])) ;
MUX2_1 m2_11 (.out(temp2[10]), .in0(temp[10]), .in1(temp[12]), .sel(dataB[1])) ;
MUX2_1 m2_12 (.out(temp2[11]), .in0(temp[11]), .in1(temp[13]), .sel(dataB[1])) ;
MUX2_1 m2_13 (.out(temp2[12]), .in0(temp[12]), .in1(temp[14]), .sel(dataB[1])) ;
MUX2_1 m2_14 (.out(temp2[13]), .in0(temp[13]), .in1(temp[15]), .sel(dataB[1])) ;
MUX2_1 m2_15 (.out(temp2[14]), .in0(temp[14]), .in1(temp[16]), .sel(dataB[1])) ;
MUX2_1 m2_16 (.out(temp2[15]), .in0(temp[15]), .in1(temp[17]), .sel(dataB[1])) ;
MUX2_1 m2_17 (.out(temp2[16]), .in0(temp[16]), .in1(temp[18]), .sel(dataB[1])) ;
MUX2_1 m2_18 (.out(temp2[17]), .in0(temp[17]), .in1(temp[19]), .sel(dataB[1])) ;
MUX2_1 m2_19 (.out(temp2[18]), .in0(temp[18]), .in1(temp[20]), .sel(dataB[1])) ;
MUX2_1 m2_20 (.out(temp2[19]), .in0(temp[19]), .in1(temp[21]), .sel(dataB[1])) ;
MUX2_1 m2_21 (.out(temp2[20]), .in0(temp[20]), .in1(temp[22]), .sel(dataB[1])) ;
MUX2_1 m2_22 (.out(temp2[21]), .in0(temp[21]), .in1(temp[23]), .sel(dataB[1])) ;
MUX2_1 m2_23 (.out(temp2[22]), .in0(temp[22]), .in1(temp[24]), .sel(dataB[1])) ;
MUX2_1 m2_24 (.out(temp2[23]), .in0(temp[23]), .in1(temp[25]), .sel(dataB[1])) ;
MUX2_1 m2_25 (.out(temp2[24]), .in0(temp[24]), .in1(temp[26]), .sel(dataB[1])) ;
MUX2_1 m2_26 (.out(temp2[25]), .in0(temp[25]), .in1(temp[27]), .sel(dataB[1])) ;
MUX2_1 m2_27 (.out(temp2[26]), .in0(temp[26]), .in1(temp[28]), .sel(dataB[1])) ;
MUX2_1 m2_28 (.out(temp2[27]), .in0(temp[27]), .in1(temp[29]), .sel(dataB[1])) ;
MUX2_1 m2_29 (.out(temp2[28]), .in0(temp[28]), .in1(temp[30]), .sel(dataB[1])) ;
MUX2_1 m2_30 (.out(temp2[29]), .in0(temp[29]), .in1(temp[31]), .sel(dataB[1])) ;
MUX2_1 m2_31 (.out(temp2[30]), .in0(temp[30]), .in1(padding), .sel(dataB[1])) ;
MUX2_1 m2_32 (.out(temp2[31]), .in0(temp[31]), .in1(padding), .sel(dataB[1])) ;

MUX2_1 m3_1 (.out(temp3[0]), .in0(temp2[0]), .in1(temp2[4]), .sel(dataB[2])) ;
MUX2_1 m3_2 (.out(temp3[1]), .in0(temp2[1]), .in1(temp2[5]), .sel(dataB[2])) ;
MUX2_1 m3_3 (.out(temp3[2]), .in0(temp2[2]), .in1(temp2[6]), .sel(dataB[2])) ;
MUX2_1 m3_4 (.out(temp3[3]), .in0(temp2[3]), .in1(temp2[7]), .sel(dataB[2])) ;
MUX2_1 m3_5 (.out(temp3[4]), .in0(temp2[4]), .in1(temp2[8]), .sel(dataB[2])) ;
MUX2_1 m3_6 (.out(temp3[5]), .in0(temp2[5]), .in1(temp2[9]), .sel(dataB[2])) ;
MUX2_1 m3_7 (.out(temp3[6]), .in0(temp2[6]), .in1(temp2[10]), .sel(dataB[2])) ;
MUX2_1 m3_8 (.out(temp3[7]), .in0(temp2[7]), .in1(temp2[11]), .sel(dataB[2])) ;
MUX2_1 m3_9 (.out(temp3[8]), .in0(temp2[8]), .in1(temp2[12]), .sel(dataB[2])) ;
MUX2_1 m3_10 (.out(temp3[9]), .in0(temp2[9]), .in1(temp2[13]), .sel(dataB[2])) ;
MUX2_1 m3_11 (.out(temp3[10]), .in0(temp2[10]), .in1(temp2[14]), .sel(dataB[2])) ;
MUX2_1 m3_12 (.out(temp3[11]), .in0(temp2[11]), .in1(temp2[15]), .sel(dataB[2])) ;
MUX2_1 m3_13 (.out(temp3[12]), .in0(temp2[12]), .in1(temp2[16]), .sel(dataB[2])) ;
MUX2_1 m3_14 (.out(temp3[13]), .in0(temp2[13]), .in1(temp2[17]), .sel(dataB[2])) ;
MUX2_1 m3_15 (.out(temp3[14]), .in0(temp2[14]), .in1(temp2[18]), .sel(dataB[2])) ;
MUX2_1 m3_16 (.out(temp3[15]), .in0(temp2[15]), .in1(temp2[19]), .sel(dataB[2])) ;
MUX2_1 m3_17 (.out(temp3[16]), .in0(temp2[16]), .in1(temp2[20]), .sel(dataB[2])) ;
MUX2_1 m3_18 (.out(temp3[17]), .in0(temp2[17]), .in1(temp2[21]), .sel(dataB[2])) ;
MUX2_1 m3_19 (.out(temp3[18]), .in0(temp2[18]), .in1(temp2[22]), .sel(dataB[2])) ;
MUX2_1 m3_20 (.out(temp3[19]), .in0(temp2[19]), .in1(temp2[23]), .sel(dataB[2])) ;
MUX2_1 m3_21 (.out(temp3[20]), .in0(temp2[20]), .in1(temp2[24]), .sel(dataB[2])) ;
MUX2_1 m3_22 (.out(temp3[21]), .in0(temp2[21]), .in1(temp2[25]), .sel(dataB[2])) ;
MUX2_1 m3_23 (.out(temp3[22]), .in0(temp2[22]), .in1(temp2[26]), .sel(dataB[2])) ;
MUX2_1 m3_24 (.out(temp3[23]), .in0(temp2[23]), .in1(temp2[27]), .sel(dataB[2])) ;
MUX2_1 m3_25 (.out(temp3[24]), .in0(temp2[24]), .in1(temp2[28]), .sel(dataB[2])) ;
MUX2_1 m3_26 (.out(temp3[25]), .in0(temp2[25]), .in1(temp2[29]), .sel(dataB[2])) ;
MUX2_1 m3_27 (.out(temp3[26]), .in0(temp2[26]), .in1(temp2[30]), .sel(dataB[2])) ;
MUX2_1 m3_28 (.out(temp3[27]), .in0(temp2[27]), .in1(temp2[31]), .sel(dataB[2])) ;
MUX2_1 m3_29 (.out(temp3[28]), .in0(temp2[28]), .in1(padding), .sel(dataB[2])) ;
MUX2_1 m3_30 (.out(temp3[29]), .in0(temp2[29]), .in1(padding), .sel(dataB[2])) ;
MUX2_1 m3_31 (.out(temp3[30]), .in0(temp2[30]), .in1(padding), .sel(dataB[2])) ;
MUX2_1 m3_32 (.out(temp3[31]), .in0(temp2[31]), .in1(padding), .sel(dataB[2])) ;

MUX2_1 m4_1 (.out(temp4[0]), .in0(temp3[0]), .in1(temp3[8]), .sel(dataB[3])) ;
MUX2_1 m4_2 (.out(temp4[1]), .in0(temp3[1]), .in1(temp3[9]), .sel(dataB[3])) ;
MUX2_1 m4_3 (.out(temp4[2]), .in0(temp3[2]), .in1(temp3[10]), .sel(dataB[3])) ;
MUX2_1 m4_4 (.out(temp4[3]), .in0(temp3[3]), .in1(temp3[11]), .sel(dataB[3])) ;
MUX2_1 m4_5 (.out(temp4[4]), .in0(temp3[4]), .in1(temp3[12]), .sel(dataB[3])) ;
MUX2_1 m4_6 (.out(temp4[5]), .in0(temp3[5]), .in1(temp3[13]), .sel(dataB[3])) ;
MUX2_1 m4_7 (.out(temp4[6]), .in0(temp3[6]), .in1(temp3[14]), .sel(dataB[3])) ;
MUX2_1 m4_8 (.out(temp4[7]), .in0(temp3[7]), .in1(temp3[15]), .sel(dataB[3])) ;
MUX2_1 m4_9 (.out(temp4[8]), .in0(temp3[8]), .in1(temp3[16]), .sel(dataB[3])) ;
MUX2_1 m4_10 (.out(temp4[9]), .in0(temp3[9]), .in1(temp3[17]), .sel(dataB[3])) ;
MUX2_1 m4_11 (.out(temp4[10]), .in0(temp3[10]), .in1(temp3[18]), .sel(dataB[3])) ;
MUX2_1 m4_12 (.out(temp4[11]), .in0(temp3[11]), .in1(temp3[19]), .sel(dataB[3])) ;
MUX2_1 m4_13 (.out(temp4[12]), .in0(temp3[12]), .in1(temp3[20]), .sel(dataB[3])) ;
MUX2_1 m4_14 (.out(temp4[13]), .in0(temp3[13]), .in1(temp3[21]), .sel(dataB[3])) ;
MUX2_1 m4_15 (.out(temp4[14]), .in0(temp3[14]), .in1(temp3[22]), .sel(dataB[3])) ;
MUX2_1 m4_16 (.out(temp4[15]), .in0(temp3[15]), .in1(temp3[23]), .sel(dataB[3])) ;
MUX2_1 m4_17 (.out(temp4[16]), .in0(temp3[16]), .in1(temp3[24]), .sel(dataB[3])) ;
MUX2_1 m4_18 (.out(temp4[17]), .in0(temp3[17]), .in1(temp3[25]), .sel(dataB[3])) ;
MUX2_1 m4_19 (.out(temp4[18]), .in0(temp3[18]), .in1(temp3[26]), .sel(dataB[3])) ;
MUX2_1 m4_20 (.out(temp4[19]), .in0(temp3[19]), .in1(temp3[27]), .sel(dataB[3])) ;
MUX2_1 m4_21 (.out(temp4[20]), .in0(temp3[20]), .in1(temp3[28]), .sel(dataB[3])) ;
MUX2_1 m4_22 (.out(temp4[21]), .in0(temp3[21]), .in1(temp3[29]), .sel(dataB[3])) ;
MUX2_1 m4_23 (.out(temp4[22]), .in0(temp3[22]), .in1(temp3[30]), .sel(dataB[3])) ;
MUX2_1 m4_24 (.out(temp4[23]), .in0(temp3[23]), .in1(temp3[31]), .sel(dataB[3])) ;
MUX2_1 m4_25 (.out(temp4[24]), .in0(temp3[24]), .in1(padding), .sel(dataB[3])) ;
MUX2_1 m4_26 (.out(temp4[25]), .in0(temp3[25]), .in1(padding), .sel(dataB[3])) ;
MUX2_1 m4_27 (.out(temp4[26]), .in0(temp3[26]), .in1(padding), .sel(dataB[3])) ;
MUX2_1 m4_28 (.out(temp4[27]), .in0(temp3[27]), .in1(padding), .sel(dataB[3])) ;
MUX2_1 m4_29 (.out(temp4[28]), .in0(temp3[28]), .in1(padding), .sel(dataB[3])) ;
MUX2_1 m4_30 (.out(temp4[29]), .in0(temp3[29]), .in1(padding), .sel(dataB[3])) ;
MUX2_1 m4_31 (.out(temp4[30]), .in0(temp3[30]), .in1(padding), .sel(dataB[3])) ;
MUX2_1 m4_32 (.out(temp4[31]), .in0(temp3[31]), .in1(padding), .sel(dataB[3])) ;

MUX2_1 m5_1 (.out(temp5[0]), .in0(temp4[0]), .in1(temp4[16]), .sel(dataB[4])) ;
MUX2_1 m5_2 (.out(temp5[1]), .in0(temp4[1]), .in1(temp4[17]), .sel(dataB[4])) ;
MUX2_1 m5_3 (.out(temp5[2]), .in0(temp4[2]), .in1(temp4[18]), .sel(dataB[4])) ;
MUX2_1 m5_4 (.out(temp5[3]), .in0(temp4[3]), .in1(temp4[19]), .sel(dataB[4])) ;
MUX2_1 m5_5 (.out(temp5[4]), .in0(temp4[4]), .in1(temp4[20]), .sel(dataB[4])) ;
MUX2_1 m5_6 (.out(temp5[5]), .in0(temp4[5]), .in1(temp4[21]), .sel(dataB[4])) ;
MUX2_1 m5_7 (.out(temp5[6]), .in0(temp4[6]), .in1(temp4[22]), .sel(dataB[4])) ;
MUX2_1 m5_8 (.out(temp5[7]), .in0(temp4[7]), .in1(temp4[23]), .sel(dataB[4])) ;
MUX2_1 m5_9 (.out(temp5[8]), .in0(temp4[8]), .in1(temp4[24]), .sel(dataB[4])) ;
MUX2_1 m5_10 (.out(temp5[9]), .in0(temp4[9]), .in1(temp4[25]), .sel(dataB[4])) ;
MUX2_1 m5_11 (.out(temp5[10]), .in0(temp4[10]), .in1(temp4[26]), .sel(dataB[4])) ;
MUX2_1 m5_12 (.out(temp5[11]), .in0(temp4[11]), .in1(temp4[27]), .sel(dataB[4])) ;
MUX2_1 m5_13 (.out(temp5[12]), .in0(temp4[12]), .in1(temp4[28]), .sel(dataB[4])) ;
MUX2_1 m5_14 (.out(temp5[13]), .in0(temp4[13]), .in1(temp4[29]), .sel(dataB[4])) ;
MUX2_1 m5_15 (.out(temp5[14]), .in0(temp4[14]), .in1(temp4[30]), .sel(dataB[4])) ;
MUX2_1 m5_16 (.out(temp5[15]), .in0(temp4[15]), .in1(temp4[31]), .sel(dataB[4])) ;
MUX2_1 m5_17 (.out(temp5[16]), .in0(temp4[16]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_18 (.out(temp5[17]), .in0(temp4[17]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_19 (.out(temp5[18]), .in0(temp4[18]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_20 (.out(temp5[19]), .in0(temp4[19]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_21 (.out(temp5[20]), .in0(temp4[20]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_22 (.out(temp5[21]), .in0(temp4[21]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_23 (.out(temp5[22]), .in0(temp4[22]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_24 (.out(temp5[23]), .in0(temp4[23]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_25 (.out(temp5[24]), .in0(temp4[24]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_26 (.out(temp5[25]), .in0(temp4[25]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_27 (.out(temp5[26]), .in0(temp4[26]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_28 (.out(temp5[27]), .in0(temp4[27]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_29 (.out(temp5[28]), .in0(temp4[28]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_30 (.out(temp5[29]), .in0(temp4[29]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_31 (.out(temp5[30]), .in0(temp4[30]), .in1(padding), .sel(dataB[4])) ;
MUX2_1 m5_32 (.out(temp5[31]), .in0(temp4[31]), .in1(padding), .sel(dataB[4])) ;

assign dataOut = ( Signal == SRL )? temp5 : 32'b0;

endmodule